`include "parallelprefix.v"
module cla16bit(a, b, Sum, cout);
    input [15:0] a, b;
    output [15:0] Sum;
    output cout;
    wire [31:0] kpg, kpg1, kpg2, kpg3, kpg4;
    wire [15:0] xor_sum, carry;
    
    assign kpg[0] = a[0];
    assign kpg[1] = b[0];
    assign kpg[2] = a[1];
    assign kpg[3] = b[1];
    assign kpg[4] = a[2];
    assign kpg[5] = b[2];
    assign kpg[6] = a[3];
    assign kpg[7] = b[3];
    assign kpg[8] = a[4];
    assign kpg[9] = b[4];
    assign kpg[10] = a[5];
    assign kpg[11] = b[5];
    assign kpg[12] = a[6];
    assign kpg[13] = b[6];
    assign kpg[14] = a[7];
    assign kpg[15] = b[7];
    assign kpg[16] = a[8];
    assign kpg[17] = b[8];
    assign kpg[18] = a[9];
    assign kpg[19] = b[9];
    assign kpg[20] = a[10];
    assign kpg[21] = b[10];
    assign kpg[22] = a[11];
    assign kpg[23] = b[11];
    assign kpg[24] = a[12];
    assign kpg[25] = b[12];
    assign kpg[26] = a[13];
    assign kpg[27] = b[13];
    assign kpg[28] = a[14];
    assign kpg[29] = b[14];
    assign kpg[30] = a[15];
    assign kpg[31] = b[15];

    assign xor_sum[0] = a[0] ^ b[0];
    assign xor_sum[1] = a[1] ^ b[1];
    assign xor_sum[2] = a[2] ^ b[2];
    assign xor_sum[3] = a[3] ^ b[3];
    assign xor_sum[4] = a[4] ^ b[4];
    assign xor_sum[5] = a[5] ^ b[5];
    assign xor_sum[6] = a[6] ^ b[6];
    assign xor_sum[7] = a[7] ^ b[7];
    assign xor_sum[8] = a[8] ^ b[8];
    assign xor_sum[9] = a[9] ^ b[9];
    assign xor_sum[10] = a[10] ^ b[10];
    assign xor_sum[11] = a[11] ^ b[11];
    assign xor_sum[12] = a[12] ^ b[12];
    assign xor_sum[13] = a[13] ^ b[13];
    assign xor_sum[14] = a[14] ^ b[14];
    assign xor_sum[15] = a[15] ^ b[15];

    parallelprefix mod0(kpg[31:30], kpg[29:28], kpg1[31:30]);
    parallelprefix mod1(kpg[29:28], kpg[27:26], kpg1[29:28]);
    parallelprefix mod2(kpg[27:26], kpg[25:24], kpg1[27:26]);
    parallelprefix mod3(kpg[25:24], kpg[23:22], kpg1[25:24]);
    parallelprefix mod4(kpg[23:22], kpg[21:20], kpg1[23:22]);
    parallelprefix mod5(kpg[21:20], kpg[19:18], kpg1[21:20]);
    parallelprefix mod6(kpg[19:18], kpg[17:16], kpg1[19:18]);
    parallelprefix mod7(kpg[17:16], kpg[15:14], kpg1[17:16]);
    parallelprefix mod8(kpg[15:14], kpg[13:12], kpg1[15:14]);
    parallelprefix mod9(kpg[13:12], kpg[11:10], kpg1[13:12]);
    parallelprefix mod10(kpg[11:10], kpg[9:8], kpg1[11:10]);
    parallelprefix mod11(kpg[9:8], kpg[7:6], kpg1[9:8]);
    parallelprefix mod12(kpg[7:6], kpg[5:4], kpg1[7:6]);
    parallelprefix mod13(kpg[5:4], kpg[3:2], kpg1[5:4]);
    parallelprefix mod14(kpg[3:2], kpg[1:0], kpg1[3:2]);
    parallelprefix mod15(kpg[1:0], 2'b00, kpg1[1:0]);

    parallelprefix mod16(kpg1[31:30], kpg1[27:26], kpg2[31:30]);
    parallelprefix mod17(kpg1[29:28], kpg1[25:24], kpg2[29:28]);
    parallelprefix mod18(kpg1[27:26], kpg1[23:22], kpg2[27:26]);
    parallelprefix mod19(kpg1[25:24], kpg1[21:20], kpg2[25:24]);
    parallelprefix mod20(kpg1[23:22], kpg1[19:18], kpg2[23:22]);
    parallelprefix mod21(kpg1[21:20], kpg1[17:16], kpg2[21:20]);
    parallelprefix mod22(kpg1[19:18], kpg1[15:14], kpg2[19:18]);
    parallelprefix mod23(kpg1[17:16], kpg1[13:12], kpg2[17:16]);
    parallelprefix mod24(kpg1[15:14], kpg1[11:10], kpg2[15:14]);
    parallelprefix mod25(kpg1[13:12], kpg1[9:8], kpg2[13:12]);
    parallelprefix mod26(kpg1[11:10], kpg1[7:6], kpg2[11:10]);
    parallelprefix mod27(kpg1[9:8], kpg1[5:4], kpg2[9:8]);
    parallelprefix mod28(kpg1[7:6], kpg1[3:2], kpg2[7:6]);
    parallelprefix mod29(kpg1[5:4], kpg1[1:0], kpg2[5:4]);
    parallelprefix mod30(kpg1[3:2], 2'b00, kpg2[3:2]);
    parallelprefix mod31(kpg1[1:0], 2'b00, kpg2[1:0]);

    parallelprefix mod32(kpg2[31:30], kpg2[23:22], kpg3[31:30]);
    parallelprefix mod33(kpg2[29:28], kpg2[21:20], kpg3[29:28]);
    parallelprefix mod34(kpg2[27:26], kpg2[19:18], kpg3[27:26]);
    parallelprefix mod35(kpg2[25:24], kpg2[17:16], kpg3[25:24]);
    parallelprefix mod36(kpg2[23:22], kpg2[15:14], kpg3[23:22]);
    parallelprefix mod37(kpg2[21:20], kpg2[13:12], kpg3[21:20]);
    parallelprefix mod38(kpg2[19:18], kpg2[11:10], kpg3[19:18]);
    parallelprefix mod39(kpg2[17:16], kpg2[9:8], kpg3[17:16]);
    parallelprefix mod40(kpg2[15:14], kpg2[7:6], kpg3[15:14]);
    parallelprefix mod41(kpg2[13:12], kpg2[5:4], kpg3[13:12]);
    parallelprefix mod42(kpg2[11:10], kpg2[3:2], kpg3[11:10]);
    parallelprefix mod43(kpg2[9:8], kpg2[1:0], kpg3[9:8]);
    parallelprefix mod44(kpg2[7:6], 2'b00, kpg3[7:6]);
    parallelprefix mod45(kpg2[5:4], 2'b00, kpg3[5:4]);
    parallelprefix mod46(kpg2[3:2], 2'b00, kpg3[3:2]);
    parallelprefix mod47(kpg2[1:0], 2'b00, kpg3[1:0]);

    parallelprefix mod48(kpg3[31:30], kpg3[15:14], kpg4[31:30]);
    parallelprefix mod49(kpg3[29:28], kpg3[13:12], kpg4[29:28]);
    parallelprefix mod50(kpg3[27:26], kpg3[11:10], kpg4[27:26]);
    parallelprefix mod51(kpg3[25:24], kpg3[9:8], kpg4[25:24]);
    parallelprefix mod52(kpg3[23:22], kpg3[7:6], kpg4[23:22]);
    parallelprefix mod53(kpg3[21:20], kpg3[5:4], kpg4[21:20]);
    parallelprefix mod54(kpg3[19:18], kpg3[3:2], kpg4[19:18]);
    parallelprefix mod55(kpg3[17:16], kpg3[1:0], kpg4[17:16]);
    parallelprefix mod56(kpg3[15:14], 2'b00, kpg4[15:14]);
    parallelprefix mod57(kpg3[13:12], 2'b00, kpg4[13:12]);
    parallelprefix mod58(kpg3[11:10], 2'b00, kpg4[11:10]);
    parallelprefix mod59(kpg3[9:8], 2'b00, kpg4[9:8]);
    parallelprefix mod60(kpg3[7:6], 2'b00, kpg4[7:6]);
    parallelprefix mod61(kpg3[5:4], 2'b00, kpg4[5:4]);
    parallelprefix mod62(kpg3[3:2], 2'b00, kpg4[3:2]);
    parallelprefix mod63(kpg3[1:0], 2'b00, kpg4[1:0]);

    assign carry[0] = kpg4[1];
    assign carry[1] = kpg4[3];
    assign carry[2] = kpg4[5];
    assign carry[3] = kpg4[7];
    assign carry[4] = kpg4[9];
    assign carry[5] = kpg4[11];
    assign carry[6] = kpg4[13];
    assign carry[7] = kpg4[15];
    assign carry[8] = kpg4[17];
    assign carry[9] = kpg4[19];
    assign carry[10] = kpg4[21];
    assign carry[11] = kpg4[23];
    assign carry[12] = kpg4[25];
    assign carry[13] = kpg4[27];
    assign carry[14] = kpg4[29];
    assign carry[15] = kpg4[31];

    assign Sum[0] = xor_sum[0];
    assign Sum[1] = xor_sum[1] ^ carry[0];
    assign Sum[2] = xor_sum[2] ^ carry[1];
    assign Sum[3] = xor_sum[3] ^ carry[2];
    assign Sum[4] = xor_sum[4] ^ carry[3];
    assign Sum[5] = xor_sum[5] ^ carry[4];
    assign Sum[6] = xor_sum[6] ^ carry[5];
    assign Sum[7] = xor_sum[7] ^ carry[6];
    assign Sum[8] = xor_sum[8] ^ carry[7];
    assign Sum[9] = xor_sum[9] ^ carry[8];
    assign Sum[10] = xor_sum[10] ^ carry[9];
    assign Sum[11] = xor_sum[11] ^ carry[10];
    assign Sum[12] = xor_sum[12] ^ carry[11];
    assign Sum[13] = xor_sum[13] ^ carry[12];
    assign Sum[14] = xor_sum[14] ^ carry[13];
    assign Sum[15] = xor_sum[15] ^ carry[14];
    assign cout = carry[15];

endmodule